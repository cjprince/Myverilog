//------------------------------------------------------------------------------------
// Copyright(c) 2022-2023 ALL rights reserved
//------------------------------------------------------------------------------------
// Author   : Lichangjiang 2452311071@qq.com
// Create   : 2023-03-10 17:14:43
// File     :  My_git_test.v
// Function : 
//------------------------------------------------------------------------------------

module My_git_test (
    
);

endmodule //My_git_test